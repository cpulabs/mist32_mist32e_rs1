// altera_asmi_rom.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module altera_asmi_rom (
		input  wire [23:0] addr,         //         addr.addr
		output wire        busy,         //         busy.busy
		input  wire        clkin,        //        clkin.clk
		output wire        data_valid,   //   data_valid.data_valid
		output wire [7:0]  dataout,      //      dataout.dataout
		input  wire        rden,         //         rden.rden
		input  wire        read,         //         read.read
		output wire [23:0] read_address, // read_address.read_address
		input  wire        reset         //        reset.reset
	);

	altera_asmi_rom_asmi_parallel_0 asmi_parallel_0 (
		.clkin        (clkin),        //        clkin.clk
		.read         (read),         //         read.read
		.rden         (rden),         //         rden.rden
		.addr         (addr),         //         addr.addr
		.reset        (reset),        //        reset.reset
		.dataout      (dataout),      //      dataout.dataout
		.busy         (busy),         //         busy.busy
		.data_valid   (data_valid),   //   data_valid.data_valid
		.read_address (read_address)  // read_address.read_address
	);

endmodule
